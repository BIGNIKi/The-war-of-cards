BIGNIK
True
77799931
